,  // ----------------------------------------------------------------------------- // Title      : I3C Slave Interface (Fully Synthesizable) // Project    : DDR5 RCD Production //----------------------------------------------------------------------------- // File       : i3c_slave_if.sv // Author     : Design Team // Revised    : 2025-11-04 // Description: Synthesizable I3C slave interface for RCD register access. //              Now supports I3C multi-beat register burst transfers (FIR/I3C burst). //              Multi-beat counting, burst handshake, packet assembly for wide mapping. //----------------------------------------------------------------------------- //////////////////////////////////////////////////////////////////////////////// // PORTS // clk, rst_n        : Clock and reset. // scl_i, sda_i      : I3C SCL/SDA inputs // scl_o, scl_oe     : SCL signal output+drive-enable (push-pull/open-drain) // sda_o, sda_oe     : SDA signal output+drive-enable (push-pull/open-drain) // static_addr       : Parameter, default static address // dynamic_addr      : Dynamic address (assigned via I3C process) // dynamic_addr_valid: Whether dynamic address is valid // current_addr      : Output, current slave address // bus_available     : True if not busy // reg_wr_en         : Pulse for register write transaction // reg_rd_en         : Pulse for register read transaction // reg_wdata         : Data to write // reg_rdata         : Data read // reg_ready         : Pulse, transaction done // rx_count/tx_count : Number of RX/TX bytes handled // err_flags         : Error status (bitfield) // burst_start       : Burst begin signal (new) // burst_end         : Burst end signal (new) // burst_beat_idx    : Beat/byte index in burst (new) // burst_size        : Burst transfer count (new) // burst_done        : Full burst done (new) // burst_ack         : Burst handshake (new) // packet_wdata      : Wide register write bus (new) // packet_rdata      : Wide register read bus (new) // packet_valid      : Packet done/valid (new) //////////////////////////////////////////////////////////////////////////////// module i3c_slave_if #(   parameter logic [6:0] STATIC_ADDR = 7'h50    
